module top;
initial begin
  $display("Hello there !!!");
  $finish;
end
endmodule
